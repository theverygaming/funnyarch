`define INITIAL_RSP 32'hFFFFFFFF
