`define INITIAL_RIP 32'hFFFFFFFF
