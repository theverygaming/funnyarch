`define INITIAL_RIP 32'h0
